library verilog;
use verilog.vl_types.all;
entity DDS_vlg_vec_tst is
end DDS_vlg_vec_tst;
